netcdf NaF_DISF {
dimensions:
	NQVALUES = 3 ;
	NTIMES = 20 ;
	NOCTANS = 8 ;
	OCTANNAME = 8 ;
	NFREQUENCIES = 20 ;
variables:
	double q(NQVALUES) ;
		q:units = "nm^-1" ;
	double time(NTIMES) ;
		time:units = "ps" ;
	char octan(NOCTANS, OCTANNAME) ;
		octan:units = "unitless" ;
	int qvectors_statistics(NQVALUES, NOCTANS) ;
	double Fqt-Na(NQVALUES, NTIMES) ;
		Fqt-Na:units = "unitless" ;
	double Fqt-total(NQVALUES, NTIMES) ;
		Fqt-total:units = "unitless" ;
	double Fqt-F(NQVALUES, NTIMES) ;
		Fqt-F:units = "unitless" ;
	double frequency(NFREQUENCIES) ;
		frequency:units = "THz" ;
	double angular_frequency(NFREQUENCIES) ;
		angular_frequency:units = "rad ps-1" ;
	double time_resolution(NFREQUENCIES) ;
		time_resolution:units = "unitless" ;
	double frequency_resolution(NFREQUENCIES) ;
		frequency_resolution:units = "unitless" ;
	double Sqw-Na(NQVALUES, NFREQUENCIES) ;
		Sqw-Na:units = "unitless" ;
	double Sqw-total(NQVALUES, NFREQUENCIES) ;
		Sqw-total:units = "unitless" ;
	double Sqw-F(NQVALUES, NFREQUENCIES) ;
		Sqw-F:units = "unitless" ;

// global attributes:
		:title = "DynamicIncoherentStructureFactor_serial" ;
		:jobinfo = "##########################################################################################\n",
			"Job information for DynamicIncoherentStructureFactor_serial analysis.\n",
			"##########################################################################################\n",
			"\n",
			"Job launched on: Mon Oct 20 17:38:50 2014\n",
			"\n",
			"General informations\n",
			"--------------------\n",
			"User: sm37\n",
			"OS: Linux-2.6.32-358.23.2.el6.x86_64\n",
			"Processor: x86_64\n",
			"nMOLDYN version: 3.0.8\n",
			"Estimate run: no\n",
			"\n",
			"Parameters\n",
			"----------\n",
			"subset = all\n",
			"timeinfo = 1:2000:100\n",
			"trajectory = /home/sm37/Projects/NaF-MD/NVT-300K/NPT-1300K/14ps/nMoldyn/NaF.nc\n",
			"qvectorsdirection = no\n",
			"pyroserver = monoprocessor\n",
			"qshellvalues = 0.0:10.0:1.0\n",
			"weights = incoherent\n",
			"deuteration = no\n",
			"qshellwidth = 1.0\n",
			"output = /home/sm37/Projects/NaF-MD/NVT-300K/NPT-1300K/14ps/nMoldyn/NaF_DISF.nc\n",
			"qvectorsgenerator = 3D isotropic\n",
			"resolution = 0.35\n",
			"qvectorspershell = 500\n",
			"\n",
			"Job status\n",
			"----------\n",
			"\n",
			"Output file written on: Mon Oct 20 17:38:50 2014\n",
			"\n",
			"" ;
data:

 q = 6, 8, 10 ;

 time = 0, 0.20000000298023224, 0.40000000596046448, 0.60000000894069672, 
    0.80000001192092896, 1.0000000149011612, 1.2000000178813934, 
    1.4000000208616257, 1.6000000238418579, 1.8000000268220901, 
    2.0000000298023224, 2.2000000327825546, 2.4000000357627869, 
    2.6000000387430191, 2.8000000417232513, 3.0000000447034836, 
    3.2000000476837158, 3.4000000506639481, 3.6000000536441803, 
    3.8000000566244125 ;

 octan =
  // octan(0, 0-7)
    "X+.Y+.Z+",
  // octan(1, 0-7)
    "X+.Y+.Z-",
  // octan(2, 0-7)
    "X+.Y-.Z+",
  // octan(3, 0-7)
    "X+.Y-.Z-",
  // octan(4, 0-7)
    "X-.Y+.Z+",
  // octan(5, 0-7)
    "X-.Y+.Z-",
  // octan(6, 0-7)
    "X-.Y-.Z+",
  // octan(7, 0-7)
    "X-.Y-.Z-" ;

 qvectors_statistics =
  // qvectors_statistics(0, 0-7)
    0, 0, 0, 1, 0, 1, 1, 3,
  // qvectors_statistics(1, 0-7)
    0, 1, 1, 2, 1, 2, 2, 3,
  // qvectors_statistics(2, 0-7)
    1, 1, 1, 1, 1, 1, 1, 1 ;

 Fqt-Na =
  // Fqt-Na(0, 0-19)
    1, 0.92811472380740201, 0.87213949738914276, 0.8212088227095754, 
    0.77783275406692887, 0.73874780735937773, 0.70916382866599792, 
    0.67897582765926445, 0.65478712865331135, 0.62709585563725945, 
    0.59626785490478906, 0.57013455260229651, 0.53121351982526122, 
    0.49980069522810933, 0.47496145484366775, 0.43954349090802203, 
    0.40648098307815206, 0.38301238199286936, 0.35496595488880472, 
    0.34597658430240363,
  // Fqt-Na(1, 0-19)
    1, 0.86210383248952782, 0.76313169241099388, 0.67847158077232794, 
    0.61283180002178494, 0.55638829370907739, 0.51065066292133254, 
    0.46692436461988313, 0.43127395201067137, 0.3969419360975785, 
    0.35358958819074782, 0.3129987177785401, 0.26337021545629369, 
    0.22880455234767227, 0.20607403447362443, 0.16802996481740126, 
    0.14017792225332162, 0.12689685437019746, 0.10351771119519099, 
    0.097069411905318481,
  // Fqt-Na(2, 0-19)
    1, 0.8014225869948256, 0.66954819425120271, 0.56468949882556729, 
    0.49243836152821624, 0.42977017364442821, 0.3778468477360955, 
    0.32713622642602125, 0.28800249113594395, 0.25586046573098115, 
    0.21389129288802194, 0.16930409260597246, 0.11657178723170304, 
    0.085853543298113899, 0.07280155905217181, 0.034439424623498902, 
    0.023615475804453209, 0.049772846283147411, 0.039598969122690703, 
    0.067676950279804193 ;

 Fqt-total =
  // Fqt-total(0, 0-19)
    0.99999999999999956, 0.92811169481436484, 0.87213269337417976, 
    0.82120025646685679, 0.7778222617959375, 0.73873188070897589, 
    0.70913949648239694, 0.67894501662638862, 0.65474777592314926, 
    0.6270496039121346, 0.59622064350233239, 0.57008342990997296, 
    0.53115886859825467, 0.49973763830696827, 0.47489214489481052, 
    0.43947931817352115, 0.40642335663781431, 0.38295336010359488, 
    0.35490898932236203, 0.34591580236687464,
  // Fqt-total(1, 0-19)
    0.99999999999999956, 0.8620983996127024, 0.7631210287479927, 
    0.67845950463752924, 0.61281769127860797, 0.55636702069777477, 
    0.51062333492213152, 0.46689108076948477, 0.43123409355993553, 
    0.39689330061213451, 0.35354001976499044, 0.31295032980668858, 
    0.26332487386721648, 0.22875417427115974, 0.20601527704114542, 
    0.16798222754636538, 0.14013743464240322, 0.12686271473703231, 
    0.10350186153380991, 0.097051061116970552,
  // Fqt-total(2, 0-19)
    0.99999999999999956, 0.80141534253317759, 0.6695361087653704, 
    0.56467737831195997, 0.49242377794911263, 0.4297494183815041, 
    0.37782540065028969, 0.32711684687927917, 0.28798277235021519, 
    0.25583411551987134, 0.21386535233532089, 0.16928428412736016, 
    0.11656510724880031, 0.085838713203058872, 0.072787279831739743, 
    0.034439663590170803, 0.023620529521296924, 0.049765967548664865, 
    0.039602880937227893, 0.067653590727241988 ;

 Fqt-F =
  // Fqt-F(0, 0-19)
    1, 0.92197798390139651, 0.85835456304418301, 0.80385361492385599, 
    0.75657541299183562, 0.70648041357393832, 0.65986682458124679, 
    0.61655267491441967, 0.5750584971678957, 0.5333898603261582, 
    0.50061755331513236, 0.46655997772479996, 0.42049013366379256, 
    0.37204737271232396, 0.3345394981465839, 0.30952953052014609, 
    0.28972981469429532, 0.26343403405684518, 0.23955371701914724, 
    0.22283238264675703,
  // Fqt-F(1, 0-19)
    1, 0.85109682401740372, 0.74152711112315306, 0.65400533161634433, 
    0.58424748628195844, 0.51328917271447538, 0.45528413641709781, 
    0.39949128356306396, 0.35052073064031702, 0.29840644236895664, 
    0.25316395738288722, 0.21496468658929466, 0.17150815578147074, 
    0.12673856910618003, 0.087031476006217925, 0.07131425348346361, 
    0.058150022350094935, 0.05772995742368324, 0.071406297165713423, 
    0.059890714629705064,
  // Fqt-F(2, 0-19)
    1, 0.78674530766400341, 0.64506299990084637, 0.54013333820298204, 
    0.46289203019897457, 0.38772001086688701, 0.33439505179711909, 
    0.28787326463944091, 0.24805223116079805, 0.20247493790383261, 
    0.16133573299884807, 0.12917211484818697, 0.10303814184071802, 
    0.055807770649816436, 0.043871858392440406, 0.034923571101879387, 
    0.033854306152642934, 0.035836530190509253, 0.047524305392726764, 
    0.02035049668345609 ;

 frequency = 0, 0.12499999813735488, 0.24999999627470976, 
    0.37499999441206461, 0.49999999254941951, 0.62499999068677436, 
    0.74999998882412922, 0.87499998696148418, 0.99999998509883903, 
    1.1249999832361939, 1.2499999813735487, 1.3749999795109036, 
    1.4999999776482584, 1.6249999757856135, 1.7499999739229684, 
    1.8749999720603232, 1.9999999701976781, 2.1249999683350329, 
    2.2499999664723878, 2.3749999646097426 ;

 angular_frequency = 0, 0.78539815169410387, 1.5707963033882077, 
    2.3561944550823113, 3.1415926067764155, 3.9269907584705188, 
    4.7123889101646226, 5.4977870618587268, 6.283185213552831, 
    7.0685833652469343, 7.8539815169410376, 8.6393796686351418, 
    9.4247778203292452, 10.21017597202335, 10.995574123717454, 
    11.780972275411557, 12.566370427105662, 13.351768578799765, 
    14.137166730493869, 14.922564882187972 ;

 time_resolution = 1, 0.99898071091997054, 0.99592907314637102, 
    0.99086371166862253, 0.98381545767196288, 0.97482703598580567, 
    0.96395263374043882, 0.9512573563244705, 0.93681657828441633, 
    0.92071519821891412, 0.90304680796896908, 0.88391278747161739, 
    0.86342133751069039, 0.84168646325244623, 0.81882692188773121, 
    0.7949651479125952, 0.7702261695670839, 0.74473652972284232, 
    0.7186232240740027, 0.69201266885627 ;

 frequency_resolution = 1, 0.0023609648579433649, 3.1071204637868238e-11, 
    2.279322120971843e-24, 9.3203530845767308e-43, 2.1244086960943744e-66, 
    2.6991239046350686e-95, 1.9115542075339542e-129, 7.5462199679007314e-169, 
    1.6605476732214969e-213, 2.0368182704994765e-263, 
    1.3926178952762632e-318, 0, 0, 0, 0, 0, 0, 0, 0 ;

 Sqw-Na =
  // Sqw-Na(0, 0-19)
    2.1496662863854685, 0.56736244022084847, 0.03436195247730111, 
    0.07664651961473154, 0.027288326627623233, 0.029857881587271973, 
    0.010242536965606621, 0.014183600016682537, 0.0083390824033198942, 
    0.0085924273358376508, 0.0056657016429464847, 0.0087479074310995442, 
    0.0024772434365405637, 0.0070691866389435646, 0.0056607554591471959, 
    0.0031380572255169433, 0.0036130087775803421, 0.0047763648545595646, 
    0.0049674370542060675, 0.0043529106994361945,
  // Sqw-Na(1, 0-19)
    1.4546884226997843, 0.6555503906440463, 0.12753236729908099, 
    0.097489053916869253, 0.063965245147499794, 0.046991319052596202, 
    0.02548787828411608, 0.024049958907575088, 0.021339909040444111, 
    0.016016183767904639, 0.010863110814089853, 0.014984052355142675, 
    0.0078295146931483383, 0.011635622084610619, 0.010758098909881194, 
    0.0064534173502319853, 0.0091594080426023877, 0.0089573375514204866, 
    0.0095348711833269303, 0.0081161558354674087,
  // Sqw-Na(2, 0-19)
    1.0642025162555124, 0.63825485173433183, 0.20381828253086623, 
    0.099745274327009831, 0.10029659779611567, 0.052094655838422217, 
    0.044248436895743322, 0.032700511141241104, 0.035351841760559423, 
    0.022915846529531898, 0.015275392106540997, 0.022354211099606319, 
    0.012645706635670821, 0.014967931589528704, 0.017204946424185113, 
    0.0073959067302346243, 0.016751540410214743, 0.01010338350573093, 
    0.016797653765451802, 0.0099515987269383731 ;

 Sqw-total =
  // Sqw-total(0, 0-19)
    2.1495417836352098, 0.56740456494072888, 0.03438157606863769, 
    0.076641923532027062, 0.027290520009762703, 0.02985458298356404, 
    0.010242582764617333, 0.014187754744433789, 0.008337917942189875, 
    0.008593327037983569, 0.0056675237531856378, 0.0087475891041923961, 
    0.0024781966860149356, 0.0070684566481143355, 0.0056602135972618319, 
    0.0031391488594492835, 0.0036129368697352584, 0.0047766077378376872, 
    0.0049668697514472105, 0.0043536869268518208,
  // Sqw-total(1, 0-19)
    1.4545819725587508, 0.65556914929653765, 0.12756296932955544, 
    0.097481736072514924, 0.06397049681736397, 0.046985507586340361, 
    0.025492710418623381, 0.024051582044986825, 0.021338713242393934, 
    0.016017651212123483, 0.010866669182844083, 0.014983261527750962, 
    0.0078309643910874725, 0.011636000875880015, 0.010756704808495927, 
    0.0064557292384691345, 0.0091577855408014434, 0.0089581131013237707, 
    0.0095345507242413797, 0.0081174932430043093,
  // Sqw-total(2, 0-19)
    1.0641575373022829, 0.63824495492156841, 0.20383374321859904, 
    0.099750804159743217, 0.10029481493086465, 0.052098457605567562, 
    0.044248556690989878, 0.032703613444571088, 0.035347224518535073, 
    0.022918566798904524, 0.015280686911340486, 0.022353253926211927, 
    0.01264654432697895, 0.014970772772899208, 0.017201886209318663, 
    0.0073993173867137304, 0.01674955344493307, 0.010105641345352048, 
    0.016794520699177681, 0.0099566926975994275 ;

 Sqw-F =
  // Sqw-F(0, 0-19)
    1.8974237138019356, 0.65270712288967114, 0.074119348613732247, 
    0.067334856035016169, 0.031732118852360852, 0.023174910460220154, 
    0.0103353257614374, 0.022601078459439972, 0.0059798841485844854, 
    0.010415223887577782, 0.0093572969958326448, 0.0081029771159374341, 
    0.0044085268758656425, 0.0055902252156367896, 0.0045629432766639859, 
    0.0053497075773264024, 0.0034673234829930479, 0.0052684463770393724, 
    0.0038180816624171182, 0.0059255474469886264,
  // Sqw-F(1, 0-19)
    1.2390204364867892, 0.69355542067702314, 0.18953208117829706, 
    0.082663101222062427, 0.074605128316077282, 0.035217288392177123, 
    0.035277782817662307, 0.027338435311001736, 0.018917222185435994, 
    0.018989225761792516, 0.018072365926296682, 0.013381836056077685, 
    0.010766602724379475, 0.012403053198288171, 0.0079336494971721794, 
    0.011137302929199646, 0.0058722193866609408, 0.010528601659054237, 
    0.0088856210745125955, 0.010825743511292228,
  // Sqw-F(2, 0-19)
    0.97307515681073697, 0.61820390903168854, 0.23514163594722182, 
    0.11094871546953894, 0.096684512789551813, 0.059797036092130586, 
    0.044491142065885537, 0.038985777701732512, 0.02599730939845632, 
    0.028427112290794185, 0.026002666654261902, 0.020414977798369406, 
    0.014342869229671033, 0.020724169111133822, 0.011004951090975663, 
    0.014305896772264796, 0.012725948740572462, 0.01467776658814412, 
    0.010450061479843935, 0.020271983309209745 ;
}
